library ieee;
use ieee.std_logic_1164.all;

package define is
  constant Enable: std_logic := '1';
  constant Disable: std_logic := '1';
  constant Zeroword: std_logic_vector := '0000000000000000';
end define;
